module top_module (input in, output out);

    not g1 (out, in);

    // assign out = !in;

endmodule